module And(
  input x,y,
  output z);

  and a1(,z,x,y);
endmodule
